// SPDX-FileCopyrightText: 2020 Efabless Corporation
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
// SPDX-License-Identifier: Apache-2.0

`default_nettype none
/*
 *-------------------------------------------------------------
 *
 * user_proj_example
 *
 * This is an example of a (trivially simple) user project,
 * showing how the user project can connect to the logic
 * analyzer, the wishbone bus, and the I/O pads.
 *
 * This project generates an integer count, which is output
 * on the user area GPIO pads (digital output only).  The
 * wishbone connection allows the project to be controlled
 * (start and stop) from the management SoC program.
 *
 * See the testbenches in directory "mprj_counter" for the
 * example programs that drive this user project.  The three
 * testbenches are "io_ports", "la_test1", and "la_test2".
 *
 *-------------------------------------------------------------
 */

module user_proj_example #(
    parameter BITS = 32,
    parameter DELAYS=10
)(
`ifdef USE_POWER_PINS
    inout vccd1,	// User area 1 1.8V supply
    inout vssd1,	// User area 1 digital ground
`endif

    // Wishbone Slave ports (WB MI A)
    input wb_clk_i,
    input wb_rst_i,
    input wbs_stb_i,
    input wbs_cyc_i,
    input wbs_we_i,
    input [3:0] wbs_sel_i,
    input [31:0] wbs_dat_i,
    input [31:0] wbs_adr_i,
    output wbs_ack_o,
    output [31:0] wbs_dat_o,

    // Logic Analyzer Signals
    input  [127:0] la_data_in,
    output [127:0] la_data_out,
    input  [127:0] la_oenb,

    // IOs
    input  [`MPRJ_IO_PADS-1:0] io_in,
    output [`MPRJ_IO_PADS-1:0] io_out,
    output [`MPRJ_IO_PADS-1:0] io_oeb,

    // IRQ
    output [2:0] irq
);
    wire clk;
    wire rst;

    wire [`MPRJ_IO_PADS-1:0] io_in;
    wire [`MPRJ_IO_PADS-1:0] io_out;
    wire [`MPRJ_IO_PADS-1:0] io_oeb;

//-----wb interface(exmem-fir)-----//
    wire valid;
    wire [3:0] wb_we;
    wire addr_decode;
    wire [(BITS-1):0] rdata;
    reg ready;
    reg [4:0] delay;//delay 10 cycle, need four bits.
//if addr = 380xxxxx, fetch instruction from user bram. 
    assign addr_decode = (wbs_adr_i[31:20] == 12'h380)? 1'b1 : 1'b0; //把wb-decode邏輯在這邊實現, 不在另外開module
    assign valid = wbs_cyc_i & wbs_stb_i & addr_decode;
    assign wb_we = wbs_sel_i & {4{wbs_we_i}};
    assign wbs_dat_o = rdata;
    assign wbs_ack_o = ready;

    always @(posedge wb_clk_i) begin
        if (wb_rst_i) begin
            ready <= 0;
            delay <= 0;
        end else begin
            ready <= 0;
            if (valid && !ready) begin
                if (delay == DELAYS - 1) begin 
                    ready <= 1;
                    delay <= 0;
                end else begin
                    delay <= delay + 1;
                end
            end
        end
    end

    bram user_bram (
        .CLK(wb_clk_i),
        .WE0(wb_we),
        .EN0(valid),
        .Di0(wbs_dat_i),
        .Do0(rdata),
        .A0(wbs_adr_i)
    );
//-----wb interface(exmem-fir)-----//


//-----wb interface(verilog fir)-----//
// implement module:WB-AXI, connect to wishbone bus signal and module:fir

//-----wb interface(verilog fir)-----//

endmodule



`default_nettype wire
